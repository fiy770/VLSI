************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: inverter_chain
* View Name:     schematic
* Netlisted on:  Oct 20 13:44:52 2016
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL	
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
*.PARAM



************************************************************************
* Library Name: VLSI
* Cell Name:    inverter
* View Name:    schematic
************************************************************************

.SUBCKT inverter1 vss vdd vin vout
*.PININFO gnd:I vdd:I vin:I vout:O
MM9 vout vin vdd vdd p_18 W=2u L=1.2u m=1 
MM8 vout vin vss vss n_18 W=0.25u L=1.2u m=1  
.ENDS
.SUBCKT inverter2 vss vdd vin vout
MM11 vout vin vdd vdd p_18 W=3.15u L=0.8u m=1 
MM10 vout vin vss vss n_18 W=0.5u L=0.8u m=1  
.ENDS
.SUBCKT inverter3 vss vdd vin vout
MM1 vout vin vdd vdd p_18 W=5u L=0.4u m=1 $8.3u 9.8u 7.1u 5.8u
MM0 vout vin vss vss n_18 W=1u L=0.4u m=1  $3u  3.5u 2.5u 2u
.ENDS
.SUBCKT inverter4 vss vdd vin vout
MM3 vout vin vdd vdd p_18 W=9.7u L=0.4u m=1 
MM2 vout vin vss vss n_18 W=2u L=0.4u m=1  
.ENDS
.SUBCKT inverter5 vss vdd vin vout
MM5 vout vin vdd vdd p_18 W=19.5u L=0.4u m=1 
MM4 vout vin vss vss n_18 W=4u L=0.4u m=1  
.ENDS
.SUBCKT inverter6 vss vdd vin vout
MM7 vout vin vdd vdd p_18 W=21.12u L=0.18u m=1 
MM6 vout vin vss vss n_18 W=8u L=0.18u m=1  
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    inverter_chain
* View Name:    schematic
************************************************************************

.SUBCKT inverter_chain vdd vin vout vss
*.PININFO vdd:I vin:I vss:I vout:O
XI1 vss vdd vin vout1  inverter1
XI2 vss vdd vout1 vout2  inverter2
XI3 vss vdd vout2 vout3  inverter3
XI4 vss vdd vout3 vout4  inverter4
XI5 vss vdd vout4 vout5  inverter5
XI6 vss vdd vout5 vout  inverter6
.ENDS

